module assert(
    input clk,
    input test
);
    always@(posedge clk)
    begin
        if(test!==1)
        begin
            $display("ASSERTION FAILED IN %m");
            $finish;
        end
    end
endmodule